//pe--pegroups-writeback
//this module is for the sum calculation and write back to the BRAM
module writeback();


endmodule