module top();




BRAMa
BRAMb

pe1 PE_(
    
);



endmodule