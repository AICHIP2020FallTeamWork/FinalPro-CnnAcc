module top();






//--------
clk_wiz_0 clk0(
);

//--------


//--------



//--------




//--------


BRAMa
BRAMb

pe1 PE(
    
);



endmodule