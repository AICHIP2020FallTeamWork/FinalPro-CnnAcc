module top(
    rst,
    clk50MHz
);


input rst;
input clk50MHz;

//-------------------------------------------

//-------------------------------------------
wire        clk;
wire        locked;
clk_wiz_0 clk0(
    .reset(rst),
    .clock_in1(clock50MHz),
    .clock_out1(clk),
    .locked(locked)
);
//-------------------------------------------




//-------------------------------------------




//-------------------------------------------





//-------------------------------------------//--------


BRAMa
BRAMb

pe1 PE(
    
);



endmodule